The leakage power of an NMOS device.

.param L = 22n
.param W = 1u
.param Vdd = 0.8
.param Vg = 0

.options noacct
.options Temp = 27

m1 d g s b nmos l={L} w={W}

vds d s {Vdd}
vgs g s {Vg}
vbs b s 0
vss s 0 0

.control
  op
  print vds#branch
.endc

.include 22nm_iHP.pm

.end
