The leakage current in a 45nm CMOS inverter.

.param Vdd = 1
.param L = 45n
.param Wp = 3u $ {4.5 * 45n}
.param Wn = 1.5u $ {1.5 * 45n}

.options Temp = 27

vdd 1 0 {Vdd}
vss 2 0 0
vin 3 0 0

x1 1 2 3 4 inv

*           vdd vss vin vout
.subckt inv 1   2   3   4
mp  pd pg ps pb pmos l={L} w={Wp}
mn  nd ng ns nb nmos l={L} w={Wn}

vpd 1  pd 0
vpg 3  pg 0
vps 4  ps 0
vpb ps pb 0

vnd 4  nd 0
vng 3  ng 0
vns 2  ns 0
vnb ns nb 0
.ends inv

.include 45nm_iHP.pm

.control
  op
  print vdd#branch
.endc

.options acct bypass=1 method=gear
.end
