The leakage power of an NMOS device.

.param L = 22n
.param W = 1u
.param Vdd = 0.8
.param Vg = 0

.options noacct
.options Temp = 27

M1 d g s b nmos l={L} w={W}

Vds d s {Vdd}
Vgs g s {Vg}
Vbs b s 0
Vss s 0 0

.control
  op
  print @M1[id]
.endc

.include 22nm_iHP.pm

.end
