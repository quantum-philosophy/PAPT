The leakage current in a CMOS inverter.

.param L = 22n
* .param Wp = {4.5 * 22n}
* .param Wn = {1.5 * 22n}
.param Wp = 2u
.param Wn = 1u

.options Temp = 27

vdd 1 0 0.8
vss 2 0 0
* vin 3 0 pulse(0 0.6 100ps 100ps 100ps 2ns 4ns)
vin 3 0 0

x1 1 2 3 4 inv

*           vdd vss vin vout
.subckt inv 1   2   3   4
mp  pd pg ps pb pmos l={L} w={Wp}
mn  nd ng ns nb nmos l={L} w={Wn}

vpd 1  pd 0
vpg 3  pg 0
vps 4  ps 0
vpb ps pb 0

vnd 4  nd 0
vng 3  ng 0
vns 2  ns 0
vnb ns nb 0
.ends inv

.include 22nm_iHP.pm

* .tran 1ps 8ns
* .op

.control
  op
  print vdd#branch
  * print vin#branch
  * print vss#branch

  * print v.x1.vnb#branch
  * print v.x1.vnd#branch
  * print v.x1.vng#branch
  * print v.x1.vns#branch

  * print @m.x1.mn[id]
  * print @m.x1.mn[ibd]
  * print @m.x1.mn[ibs]
  * print @m.x1.mn[isub]
  * print @m.x1.mn[igs]
  * print @m.x1.mn[igd]
  * print @m.x1.mn[igb]
  * print @m.x1.mn[igcs]
  * print @m.x1.mn[igcd]

  * print v.x1.vpb#branch
  * print v.x1.vpd#branch
  * print v.x1.vpg#branch
  * print v.x1.vps#branch

  * print @m.x1.mp[id]
  * print @m.x1.mp[ibd]
  * print @m.x1.mp[ibs]
  * print @m.x1.mp[isub]
  * print @m.x1.mp[igs]
  * print @m.x1.mp[igd]
  * print @m.x1.mp[igb]
  * print @m.x1.mp[igcs]
  * print @m.x1.mp[igcd]
.endc

.options acct bypass=1 method=gear
.end
